context work.test_contaext;
library IEEE;
context IEEE.IEEE_STD_CONTEXT;
entity test is
end entity;