entity ent is
  port (
    apple: inout integer -- vhdl-linter-disable-line unused
  );
end entity;
architecture arch of ent is
begin
end architecture;