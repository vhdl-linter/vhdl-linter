use work.util.all;

entity ent is
  !declaration
end;