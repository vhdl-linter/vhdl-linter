
entity ent is
end;
architecture rtl of ent is
  procedure p;
begin
  !statement
end;
