entity test is
end entity;
architecture rtl of test is

begin
end architecture; 