entity ent is
end entity;
architecture arch of ent is
  signal apple: integer; -- vhdl-linter-disable-line unused
begin
end architecture;