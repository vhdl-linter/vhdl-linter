library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ent is
  port (
    o_test : out unsigned(1 downto 0)
    );
end ent;
