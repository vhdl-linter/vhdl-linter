entity foo is
end entity;
