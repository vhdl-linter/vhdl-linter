context test_contextA is
  library test_03_library;

  context test_03_library.test_ContextB;
end context;