entity test is
  port (
    );
end test;
architecture arch of test is
begin
  p_gen : if true generate

  else generate

  end generate;
end arch;
