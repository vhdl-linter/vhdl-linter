entity sub is
end entity;
architecture rtl of sub is
begin
end architecture;