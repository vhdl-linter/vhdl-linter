entity ent is
end entity;
architecture arch of ent is
  signal apple: integer;
begin
end architecture;