library ieee;

package pkg is
  use ieee; -- expect a package
end package;