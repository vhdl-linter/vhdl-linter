library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
entity test_use is
end entity;
architecture arch of test_use is
  signal a : std_ulogic;
begin
end architecture;
