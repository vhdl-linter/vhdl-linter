
context test_contextB is
  library test_02_deallocate;
  use test_02_deallocate.deallocate_test_pkg_def.all;
end context;
