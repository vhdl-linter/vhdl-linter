
entity architecture_begin_missing is

end architecture_begin_missing ;

architecture arch of architecture_begin_missing is

-- begin
  assert true report "ASD";
end architecture ;