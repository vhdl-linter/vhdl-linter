-- Based on #178

library ieee;
use ieee.std_logic_1164.all;

entity test_arch is
end entity;
architecture arch of test_arch is

begin
  foo <= '01';
end arch;
