library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_entity is
end test_entity;

architecture arch of test_entity is

begin
end architecture arch;
