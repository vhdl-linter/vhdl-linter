entity test is
end test;
architecture arch of test is
  --vhdl-linter-disable-next-line unused
  signal test : integer;

begin
test <= 0;
end arch ;