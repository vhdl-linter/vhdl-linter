entity exit is -- exit is reserved word/keyword
end exit;