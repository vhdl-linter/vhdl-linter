package deallocate_test_pkg_def is
  type test_type is access integer;

end package;
