context test_contextA is
  library test_deallocate;

  context test_deallocate.test_contextB;
end context;
