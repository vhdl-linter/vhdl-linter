-- Dummy for other test cases.
entity test is
  port (
    i : in std_logic -- dummy error
  );
end entity;
context test_ContextB is
end context;