library test_03_library;
use test_03_library.foo.all;
entity test is
end entity;
