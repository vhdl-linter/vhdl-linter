context work.contextA;
entity dummy is
end entity;


architecture arch of dummy is
  constant TEST_VAR : integer := TEST_CONSTANT + 1;
begin

end architecture;
