architecture arch of units is -- units is reserved
begin
  a_p : process
  begin
    wait for 6 ns;
  end process;
end architecture;
