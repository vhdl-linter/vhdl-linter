context test_contextA is
  context work.test_ContextB;
end context;
