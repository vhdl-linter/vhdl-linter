entity test_inst1 is
end entity;
architecture r of test_inst1 is
begin
 i: entity work.test_vhdl;
end architecture;