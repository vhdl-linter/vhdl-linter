library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ent is

end ent;

architecture arch of ent is



  attribute PIN_NO unexpected;

begin

end architecture;

entity adder is
end entity;
