entity test_tool_reporting is
end entity;
architecture arch of test_tool_reporting is
begin
  `warning "yoyoyo"
end architecture;