package dummy_pkg is
  constant a : NOT_EXIST; -- dummy error
end package;