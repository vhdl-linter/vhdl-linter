entity ent is
  port (
    apple: in integer
  );
end entity;
architecture arch of ent is
begin
end architecture;