-- library test;
use test.foo.all;
entity test_entity is
end entity;
