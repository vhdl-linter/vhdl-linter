library test_lib;

entity test2 is
end entity;

architecture arch of test2 is


begin
  inst_test : entity test_lib.test;

end;
