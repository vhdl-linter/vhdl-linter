entity test_inst is
end entity;
architecture rtl of test_inst is
begin
  inst: entity work.test_entity_b;
end architecture;