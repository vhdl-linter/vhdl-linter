architecture arch of asd  is


begin

end arch;
