package pkg is
  constant apple: integer := 2;
end;