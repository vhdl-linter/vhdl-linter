library ieee;
use ieee.std_logic_1164.all;

entity ent is
end ent;
architecture arch of ent is

  signal test_unused : std_ulogic;

begin

end arch ; -- arch
