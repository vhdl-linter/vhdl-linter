

entity test_inst is
end test_inst;

architecture arch of test_inst is
begin
  test_inst : entity work.test_entity;
end architecture;
