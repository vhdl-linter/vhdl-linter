entity test_inst2 is
end entity;
architecture r of test_inst2 is
begin
 i: entity work.test_verilog;
end architecture;