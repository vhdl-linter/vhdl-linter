context test_contextA is
  context test.test_ContextB;
end context;
