entity test_entity_a is
end entity;