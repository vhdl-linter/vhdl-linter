package pkg is
  constant a : integer := 5;

pkg;



package body pkg is

pkg;

package pkg2 is
  constant a : integer := 5;
;
package body pkg2 is
;
