use work.util.all;

entity ent is
end;
architecture rtl of ent is
begin
  process
    !declaration
  begin
  end process;
end;