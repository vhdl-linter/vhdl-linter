entity ent is
  generic (
    apple: integer
  );
end entity;
architecture arch of ent is
begin
end architecture;