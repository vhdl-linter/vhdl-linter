entity empty_interface_list_parameter is
  procedure dummy ()
  is
  begin
  end procedure;
begin
end entity;
