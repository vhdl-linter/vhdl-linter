entity torture_entity is
end torture_entity;

architecture arch of torture_entity is
signal a : integer;
signal b : integer;
begin
    a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;
  a <= b;

end architecture;
