library ieee;
context ieee.ieee_std_context;
entity test_context is
end entity;
architecture arch of test_context is
  signal a : std_ulogic;
begin
end architecture;
