library ieee, test;
use ieee.std_logic_1164.all;
use std.textio.all;

entity test_library_list is
end entity;
architecture arch of test_library_list is
begin
end architecture;
