library ieee;
use ieee.std_logic_1164.all;

entity ent is
  port (
    o_test : out std_ulogic_vector(1 downto 0)
    );
end ent;
