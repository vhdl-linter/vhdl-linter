package test_pkg is

end package test_pkg;
package body test_pkg is
end package body test_pkg;
