--vhdl-linter-disable multiple-definition
entity ignore_file is
  port (
    input : integer
    );
end entity;
architecture rtl of ignore_file is
begin

end architecture;
