library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pkg is
  function func(
    a: integer;
    b: integer
  ) return integer;
end package;  