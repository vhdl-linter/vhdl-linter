entity semicolon_generic_list is
  generic (
    input : std_logic;
    );
end entity;
