library ieee;
use ieee.std_logic_1164.all;
entity test_entity is
  port (
    clk_in : std_ulogic
    );
end entity;
