--! @library libA
package test_package is
end package;