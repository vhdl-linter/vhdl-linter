entity test_use is
end entity;
architecture arch of test_use is
begin
  inst: entity work.test_entity;
end architecture;