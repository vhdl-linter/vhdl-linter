context test_contextA is
  library test;

  context test.test_ContextB;
end context;
