--! @library libA
entity test_entity is
end test_entity;
configuration test_entity_cfg of test_entity is
end configuration;