entity test_entity_b is
end entity;