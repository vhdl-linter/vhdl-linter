entity semicolon_parameter_list is
  procedure dummy parameter -- If parameter keyword is used there need to be a parameter list
  is
  begin
  end procedure;
begin
end entity;
