library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pkg_test_inner is

  type test_record_inner is record
    foo_inner : integer;
  end record;
  type test_record is record
    foo : test_record_inner;
  end record;

end package;
