context test_contextA is
  library test_02_deallocate;

  context test_02_deallocate.test_ContextB;
end context;
