package pkg is
  procedure proc(
    apple: out integer -- vhdl-linter-disable-line unused
  );
end package;