library ieee;

entity ent is

  use ieee.numeric_std.all;

end entity;