
context test_contextB is
  library test_deallocate;
  use test_deallocate.deallocate_test_pkg_def.all;
end context;
