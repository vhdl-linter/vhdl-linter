entity test is
end entity;
architecture arch of test is
begin
end architecture;