
      module test_enttity
      endmodule;