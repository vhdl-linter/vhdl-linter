library test_library;
use test_library.foo.all;
entity test is
end entity;
