library ieee;
use ieee.std_logic_1164.all;
entity info is
  port (
    apple: in std_logic -- resolved
  );
end entity;