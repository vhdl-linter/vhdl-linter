
entity test_entity_split is
  port (
    foo : in integer
    );
end test_entity_split;
