package error is
  constant s : std_ulogic := '2'; -- std_ulogic not imported
end package;
