module test_multiple_module1
#(
  parameter WIDTH = 8
)
(
		input  wire [0:0]   in_bit,
		output wire [0:0]   out_bit // test comment
    );
endmodule;
module test_multiple_module2
#(
  parameter WIDTH = 8
)
(
		input  wire [0:0]   in_bit2,
		output wire [0:0]   out_bit2 // test comment
    );
endmodule;