entity units is
end units ;

architecture arch of units is

begin
  a_p: process
  begin
        wait for 6 ns ;
end process;

end architecture ;