-- library test;
use test.foo.all;
entity test is
end entity;
