entity ent is
end entity;
architecture arch of ent is
begin
  apple: entity work.ent;
end architecture;