use work.util.all;

package pkg is
end package;
package body pkg is
  procedure x is
    !declaration
  begin
  end procedure;
end ;