
      entity test_entity is
      end entity;