entity test is
  port (

  );
end entity;
architecture arch of test is
begin
end architecture;