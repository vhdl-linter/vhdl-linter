entity test_vhdl is
end entity;
architecture rtl of test_vhdl is
begin
 -- this is a long comment to make the file too large
 -- Lorem ipsum dolor sit amet, consectetur adipiscing elit. Etiam ipsum mauris, consectetur nec nisl id, finibus commodo sem. Phasellus eu quam blandit, pulvinar metus sed, suscipit elit. Donec porta, lacus vel elementum elementum, elit sem tempus eros, a commodo massa metus id elit. Etiam tristique commodo urna, ut malesuada tortor malesuada facilisis. Phasellus ultricies, lectus ut accumsan congue, massa sapien iaculis nunc, id porttitor purus justo sed massa. Sed posuere purus massa, sed gravida erat faucibus eget. Suspendisse porta dui ac leo sodales euismod. In scelerisque dui quis faucibus malesuada. Duis a rhoncus erat. Nam id viverra sem, et pretium velit. Quisque dignissim, erat eget dapibus ullamcorper, mi sem eleifend turpis, sit amet iaculis turpis diam vitae erat. Donec pellentesque luctus malesuada. Vestibulum vulputate nunc sit amet enim pretium posuere. Donec ultrices mauris vitae volutpat tristique. Nunc dui augue, fringilla a commodo id, tristique et ipsum. 
end architecture;