package pkg is
  procedure proc(
    apple: inout integer -- vhdl-linter-disable-line unused
  );
end package;