entity warning is
  port (
    input: in integer -- unused
  );
end entity;
architecture rtl of warning is
begin
end architecture;