entity ignore_line is
  port (
    input : integer  --vhdl-linter-disable-line multiple-definition
    );
end entity;
architecture rtl of ignore_line is
begin

end architecture;
