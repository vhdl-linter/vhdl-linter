entity dummy is

end dummy;
architecture arch of dummy is

  signal a_unused : std_ulogic;

begin

end arch ; -- arch