
context test_contextB is
  library test_lib;
  use test_lib.deallocate_test_pkg_def.all;
end context;
