context work.test_context;
entity use_context is
end entity;
architecture arch of use_context is
  signal a : t_enum;
begin

end architecture;
