
context test_contextB is
  use work.deallocate_test_pkg_def.all;
end context;
