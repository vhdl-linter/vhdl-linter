--vhdl-linter-disable
entity test is
end test;
architecture arch of test is
  signal test : integer;

begin
  test <= 0;
end arch;
