context test_context is
  use work.test_pkg.all;
end context test_context;