entity test is
end test;
architecture arch of test is
  signal test : integer; --vhdl-linter-disable-line unused

begin
test <= 0;
end arch ;