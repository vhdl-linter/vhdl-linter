
entity port_integer_range is
  port (
    i_i: in integer range 0 to 10
  );
end entity;

