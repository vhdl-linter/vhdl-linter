context test_context is
  use work.deallocate_test_pkg_def.all;
end context;
