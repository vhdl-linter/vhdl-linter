entity test_hover is
  `if VALUE5 > "5" then
    `error "FALSE"
  `end if
end entity;