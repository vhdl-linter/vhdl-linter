use work.util.all;

package pkg is
  type t is protected
  end protected;
end package;
package body pkg is
  type t is protected body
    !declaration
  end protected body;
end package body;