
entity test_entity_split is
end test_entity_split ;