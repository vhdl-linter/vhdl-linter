package pkg is
  variable apple: integer;
end;