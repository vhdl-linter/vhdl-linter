library IEEE;
use work.util.all;

configuration conf of xyz is
  !declaration
end configuration;
