-- vhdl-linter-disable port-declaration
entity pkg_in_port_map is
end entity;
architecture arch of pkg_in_port_map is
  subtype test_unused is work.dummy_pkg;
begin

end architecture;
