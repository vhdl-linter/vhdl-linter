entity ent is
procedure p;
begin
  !statement
end;