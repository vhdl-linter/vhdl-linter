entity component_entity is
  port(
    i_clk: in integer
  );
end entity component_entity;