
package instantiated_pkg is new work.generic_pkg; 