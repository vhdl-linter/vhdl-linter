package test is
  alias SIGN : bit is bit_vector(0 to 31);
  alias test is sign;
end package;
