
context test_contextB is
  library test;
  use test.deallocate_test_pkg_def.all;
end context;
