
context test_contextB is
  use test.deallocate_test_pkg_def.all;
end context;
