package foo is
  constant a : integer; -- dummy error
end package;
context test_contextB is
end context;