package test_pkg is

end package;