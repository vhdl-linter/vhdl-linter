context test_contextA is
  library test_lib;

  context test.test_ContextB;
end context;
