entity entity_name is

end entity;
architecture arch of does_not_exist is -- entity name wrong, will not find entity
begin
end architecture;
