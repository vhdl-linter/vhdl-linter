library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_completion is

end test_completion;

architecture arch of test_completion is
  signal a : STD_LOGIC;
begin

end arch;
