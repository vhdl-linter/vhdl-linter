entity test is
end entity;
architecture arch of test is
  use work.test_pkg.all; -- test_pkg does not exist

begin
end arch;