entity ent is
  port (
    apple: inout integer
  );
end entity;
architecture arch of ent is
begin
end architecture;