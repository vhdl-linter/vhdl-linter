package pkg is
  procedure proc(
    apple: in integer -- vhdl-linter-disable-line unused
  );
end package;