entity empty_interface_list is
  port ( -- Empty interface list
  );
end entity;
