entity test_instantiation is
end entity;
architecture arch of test_instantiation is
begin
test_entity : entity work.test_entity;

end architecture;