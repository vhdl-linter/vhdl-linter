context test_contextA is
  library test_library;

  context test_library.test_contextB;
end context;