library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_alias_procedure is
end test_alias_procedure;

architecture arch of test_alias_procedure is

  alias test_alias is ; -- name is missing
begin

end architecture;
