entity generic_entity is
  generic (
    GENERIC_NAME : integer
  );
end generic_entity;