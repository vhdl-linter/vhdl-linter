entity ent is
  port (
    apple: out integer
  );
end entity;
architecture arch of ent is
begin
end architecture;