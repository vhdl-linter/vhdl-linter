package protected_Type is

end package;
package body protected_Type is


end package body;