library ieee;
use ieee.std_logic_1164.all;
entity attribute_missing_prefix is

end entity;
architecture arch of attribute_missing_prefix is
  -- signal b : slv_vector(range a'range);
  -- signal b : std_ulogic_vector(a');
begin
end architecture;
