�.����+r�#9�˂��8�$0�����7O&���*�]o�^�l:h���0\�uP��OW�����^�,���鳋Nc�+�A��7:kB�"�����@��]h�>��Hv���2Sqnf����V@[�0�&"PF���]gr0H$3��RJ�Z�L��[���..�e��C�{�����ǅ�Ǝ�a�~
��Μ����0"mlC�(T�'X��AfK	�f��
��L�DAD�d��~1����5O:�SX���=Y����2~Qd!���ػ��C��5�Ɔ��0Ǘh����
y�� �Vx��s�n��QE��/��m�+���%�4�0�*x�'V��;Է�E���R��~���C=�%P�y/�|�[�?�5���FWw��9y�' ���3@��p�G%W�J�����21䋫����|ؐS^�7ICLZU�����)��2^Wڔ��yJ"f���� >�3PEM4�� '���"Y��t%�F�r%v�4��=Ms��R�+����?���Y�k���U�HW3D�,�m��Տ�Y6S���97�)��f57uT��N����EF��
�:��] $��Qm^�!;deA�̱ڬ5T`ek�x���J,:�@%1��҂s�*��Q�7Y�%���4���G�G�	��UL�@�B��P�LeX
=r�{UM;�����ul��9�T�������A���BYj'�d��E��T6(��]�����0}^ظ���o�"q��CD|�$mq�5�,@;ȭ5��Ǽ�k#�ALkT ��D6�X�a �x� e����$˶�0,̓�<�-Д���HN4��*Ի�����2�)��g��6�	 �oqO��K�� rW@�i9�7m��L�	��|���!pk��S�+�{����'pR@4$rJ�$�.畻׍�U��"�F(A����M��N��q����^����ہ��Ė$�)Ż��En�� i徕jlMJn�HB� �m