library ieee;
use ieee.std_logic_1164.all;

package pkg is
  type x is record
    child: std_ulogic;
  end record;
end package;
