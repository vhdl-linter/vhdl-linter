library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pkg_test is
  constant a : no_exists; -- dummy error
end package;