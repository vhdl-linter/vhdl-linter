library ieee;
entity dummy is
end dummy;
architecture arch of dummy is

begin
  p_test : process
  begin
    report CopyRightNotice;
  end process;
end arch;  -- arch
