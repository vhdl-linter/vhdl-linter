use work.util.all;

package pkg is
  !declaration
end package;