entity test_entity is

end test_entity;