entity test_entity is
  generic (
    i_a : in integer
    );

end entity;
