entity empty_interface_list_generic is
  generic ( -- Empty interface list
  );
end entity;
