-- File contains only comment