package error is
  constant s : std_ulogic := '1'; -- std_ulogic not imported
end package;
