use work.util.all;

package pkg is
end package;
package body pkg is
  !declaration
end ;