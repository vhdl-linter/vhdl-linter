library IEEE;
entity dummy is
  port (
    i_foo : std_ulogic
    );
end dummy;
