-- vhdl-linter-disable port-declaration
library ieee;
use ieee.std_logic_1164.NOT_EXIST; --is not part of the package
entity test_not_all is
end test_not_all;
