package foo is
  constant a : integer; -- dummy error
end package;
