package foo is
  constant a : no_exists; -- dummy error
end package;
