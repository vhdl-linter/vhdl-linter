architecture arch of test_entity_split  is


begin

end arch;
