package body pkg_no_header is
end package body;