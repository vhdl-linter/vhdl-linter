-- Test case for fixed bug where a broken vhdl file in the same folder broke the renaming logic
use std.textio.all;
use work.stop_pkg;
package dummy is
end package;