use work.util.all;

package pkg is
  type t is protected
    !declaration
  end protected;
end package;