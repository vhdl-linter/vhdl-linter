package generic_pkg is
  generic (
    generic_parameter : integer := 0
    ) --dummy error
end package;