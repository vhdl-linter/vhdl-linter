library ieee;
use ieee.std_logic_1164.all;
entity foo is
  port (
    i_a : out std_ulogic
    );
end entity;