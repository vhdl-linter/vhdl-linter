context test_contextA is
  library test_lib;

  context test_lib.test_ContextB;
end context;
