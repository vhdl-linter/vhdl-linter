
architecture arch of foo is
begin
  apple.kiwi;
end arch;
