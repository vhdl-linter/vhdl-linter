library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
entity test_line is
end entity;
architecture arch of test_line is

  alias BREAD is READ [line, std_ulogic_vector, boolean, STD_ULOGIC];

begin
end architecture;
