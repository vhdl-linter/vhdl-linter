library ieee;
use ieee.std_logic_1164.all;
entity type_in_interface_pkg is
generic (
  package test_pkg is new std_ulogic generic map (<>)
  );

end entity;