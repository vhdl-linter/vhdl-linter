configuration dut_cfg of for_test is
  for arch
  end for;
end configuration;