

package pkg is
  -- package inner is
  -- end package;
end package;