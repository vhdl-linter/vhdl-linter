-- test_04_generic_package
package instantiated_pkg is new test_04_generic_package.generic_pkg;