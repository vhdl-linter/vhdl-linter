entity semicolon_port_list is
  port (
    input : in std_logic;
    );
end entity;
