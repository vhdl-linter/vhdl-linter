use work.util.all;

entity ent is
end;
architecture rtl of ent is
  !declaration
begin
end;