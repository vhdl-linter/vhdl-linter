-- Dummy for other test cases.
entity test is
  port (
    i_a : in std_ulogic -- dummy error
  );
end entity;
context test_ContextB is
end context;