context recursive_context is
  library ieee;
  context ieee.ieee_std_context;
end context;
