entity port_range_2 is
  port (
    i_i: in integer range 0 to integer'high
  );
end entity;