-- placeholder entity
entity foo is
end entity;