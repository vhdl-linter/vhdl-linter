architecture arch of test_entity_split  is
 signal bar : integer;

begin
  bar <= foo;
end arch;
