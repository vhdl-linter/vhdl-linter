entity test is
end entity;
architecture arch of test is
  use work.test_pkg.all; -- work. should not be here

begin
end arch;